package psw_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "seq_trans.sv"
`include "config_psw.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agt.sv"
`include "sequence_base.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"
endpackage::psw_pkg